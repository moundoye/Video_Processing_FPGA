// elimax_ghrd_nios_sys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module elimax_ghrd_nios_sys (
		input  wire        altpll_0_areset_conduit_export,                       //                altpll_0_areset_conduit.export
		output wire        altpll_0_c0_clk,                                      //                            altpll_0_c0.clk
		output wire        altpll_0_locked_conduit_export,                       //                altpll_0_locked_conduit.export
		output wire        clear_external_connection_export,                     //              clear_external_connection.export
		input  wire        clk_clk,                                              //                                    clk.clk
		output wire        clock_bridge_0_out_clk_clk,                           //                 clock_bridge_0_out_clk.clk
		output wire [1:0]  led_external_connection_export,                       //                led_external_connection.export
		inout  wire        opencores_i2c_0_export_0_scl_pad_io,                  //               opencores_i2c_0_export_0.scl_pad_io
		inout  wire        opencores_i2c_0_export_0_sda_pad_io,                  //                                       .sda_pad_io
		input  wire        reset_reset_n,                                        //                                  reset.reset_n
		output wire        trigger_external_connection_export,                   //            trigger_external_connection.export
		input  wire [7:0]  usb_streaming_0_asi_in0_data,                         //                usb_streaming_0_asi_in0.data
		input  wire        usb_streaming_0_asi_in0_endofpacket,                  //                                       .endofpacket
		input  wire        usb_streaming_0_asi_in0_startofpacket,                //                                       .startofpacket
		input  wire        usb_streaming_0_asi_in0_valid,                        //                                       .valid
		input  wire        usb_streaming_0_clear_fifo_conduit,                   //             usb_streaming_0_clear_fifo.conduit
		output wire        usb_streaming_0_ctl0_conduit,                         //                   usb_streaming_0_ctl0.conduit
		output wire        usb_streaming_0_ctl1_conduit,                         //                   usb_streaming_0_ctl1.conduit
		output wire        usb_streaming_0_ctl11_conduit,                        //                  usb_streaming_0_ctl11.conduit
		output wire        usb_streaming_0_ctl12_conduit,                        //                  usb_streaming_0_ctl12.conduit
		output wire        usb_streaming_0_ctl2_conduit,                         //                   usb_streaming_0_ctl2.conduit
		output wire        usb_streaming_0_ctl3_conduit,                         //                   usb_streaming_0_ctl3.conduit
		input  wire        usb_streaming_0_ctl4_sw_conduit,                      //                usb_streaming_0_ctl4_sw.conduit
		input  wire        usb_streaming_0_ctl5_conduit,                         //                   usb_streaming_0_ctl5.conduit
		input  wire        usb_streaming_0_ctl6_conduit,                         //                   usb_streaming_0_ctl6.conduit
		output wire        usb_streaming_0_ctl7_conduit,                         //                   usb_streaming_0_ctl7.conduit
		input  wire        usb_streaming_0_ctl8_conduit,                         //                   usb_streaming_0_ctl8.conduit
		inout  wire [15:0] usb_streaming_0_usb_data_conduit,                     //               usb_streaming_0_usb_data.conduit
		input  wire [3:0]  usbstatus_external_connection_export,                 //          usbstatus_external_connection.export
		output wire [7:0]  videosampler_0_avalon_streaming_source_data,          // videosampler_0_avalon_streaming_source.data
		output wire        videosampler_0_avalon_streaming_source_valid,         //                                       .valid
		output wire        videosampler_0_avalon_streaming_source_endofpacket,   //                                       .endofpacket
		output wire        videosampler_0_avalon_streaming_source_startofpacket, //                                       .startofpacket
		input  wire        videosampler_0_href_conduit,                          //                    videosampler_0_href.conduit
		input  wire        videosampler_0_pclk_i_conduit,                        //                  videosampler_0_pclk_i.conduit
		input  wire [7:0]  videosampler_0_pixel_i_conduit,                       //                 videosampler_0_pixel_i.conduit
		input  wire        videosampler_0_vsync_i_conduit                        //                 videosampler_0_vsync_i.conduit
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                            // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                         // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [18:0] nios2_gen2_0_data_master_address;                             // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                          // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                               // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                           // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [18:0] nios2_gen2_0_instruction_master_address;                      // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                         // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect;  // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_chipselect -> opencores_i2c_0:wb_stb_i
	wire   [7:0] mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata;    // opencores_i2c_0:wb_dat_o -> mm_interconnect_0:opencores_i2c_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_opencores_i2c_0_avalon_slave_0_waitrequest; // opencores_i2c_0:wb_ack_o -> mm_interconnect_0:opencores_i2c_0_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address;     // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_address -> opencores_i2c_0:wb_adr_i
	wire         mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write;       // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_write -> opencores_i2c_0:wb_we_i
	wire   [7:0] mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata;   // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_writedata -> opencores_i2c_0:wb_dat_i
	wire  [31:0] mm_interconnect_0_videosampler_0_avalon_slave_0_readdata;     // videosampler_0:datard_o -> mm_interconnect_0:videosampler_0_avalon_slave_0_readdata
	wire   [2:0] mm_interconnect_0_videosampler_0_avalon_slave_0_address;      // mm_interconnect_0:videosampler_0_avalon_slave_0_address -> videosampler_0:addr_rel_i
	wire         mm_interconnect_0_videosampler_0_avalon_slave_0_read;         // mm_interconnect_0:videosampler_0_avalon_slave_0_read -> videosampler_0:rd_i
	wire         mm_interconnect_0_videosampler_0_avalon_slave_0_write;        // mm_interconnect_0:videosampler_0_avalon_slave_0_write -> videosampler_0:wr_i
	wire  [31:0] mm_interconnect_0_videosampler_0_avalon_slave_0_writedata;    // mm_interconnect_0:videosampler_0_avalon_slave_0_writedata -> videosampler_0:datawr_i
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;        // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;         // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;      // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;   // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;          // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                 // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                    // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                   // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;               // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_trigger_s1_chipselect;                      // mm_interconnect_0:trigger_s1_chipselect -> trigger:chipselect
	wire  [31:0] mm_interconnect_0_trigger_s1_readdata;                        // trigger:readdata -> mm_interconnect_0:trigger_s1_readdata
	wire   [2:0] mm_interconnect_0_trigger_s1_address;                         // mm_interconnect_0:trigger_s1_address -> trigger:address
	wire         mm_interconnect_0_trigger_s1_write;                           // mm_interconnect_0:trigger_s1_write -> trigger:write_n
	wire  [31:0] mm_interconnect_0_trigger_s1_writedata;                       // mm_interconnect_0:trigger_s1_writedata -> trigger:writedata
	wire         mm_interconnect_0_clear_s1_chipselect;                        // mm_interconnect_0:clear_s1_chipselect -> clear:chipselect
	wire  [31:0] mm_interconnect_0_clear_s1_readdata;                          // clear:readdata -> mm_interconnect_0:clear_s1_readdata
	wire   [1:0] mm_interconnect_0_clear_s1_address;                           // mm_interconnect_0:clear_s1_address -> clear:address
	wire         mm_interconnect_0_clear_s1_write;                             // mm_interconnect_0:clear_s1_write -> clear:write_n
	wire  [31:0] mm_interconnect_0_clear_s1_writedata;                         // mm_interconnect_0:clear_s1_writedata -> clear:writedata
	wire         mm_interconnect_0_led_s1_chipselect;                          // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                            // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                             // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                               // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                           // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_usbstatus_s1_chipselect;                    // mm_interconnect_0:usbstatus_s1_chipselect -> usbstatus:chipselect
	wire  [31:0] mm_interconnect_0_usbstatus_s1_readdata;                      // usbstatus:readdata -> mm_interconnect_0:usbstatus_s1_readdata
	wire   [1:0] mm_interconnect_0_usbstatus_s1_address;                       // mm_interconnect_0:usbstatus_s1_address -> usbstatus:address
	wire         mm_interconnect_0_usbstatus_s1_write;                         // mm_interconnect_0:usbstatus_s1_write -> usbstatus:write_n
	wire  [31:0] mm_interconnect_0_usbstatus_s1_writedata;                     // mm_interconnect_0:usbstatus_s1_writedata -> usbstatus:writedata
	wire         irq_mapper_receiver0_irq;                                     // opencores_i2c_0:wb_inta_o -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                         // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [clear:reset_n, jtag_uart_0:rst_n, led:reset_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, opencores_i2c_0:wb_rst_i, rst_translator:in_reset, sysid_qsys_0:reset_n, trigger:reset_n, usb_streaming_0:reset_n, usbstatus:reset_n, videosampler_0:reset_n_i]
	wire         rst_controller_001_reset_out_reset_req;                       // rst_controller_001:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                           // rst_controller_002:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                       // rst_controller_002:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                       // nios2_gen2_0:debug_reset_request -> rst_controller_002:reset_in1

	elimax_ghrd_nios_sys_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.c1                 (clock_bridge_0_out_clk_clk),                     //                    c1.clk
		.areset             (altpll_0_areset_conduit_export),                 //        areset_conduit.export
		.locked             (altpll_0_locked_conduit_export),                 //        locked_conduit.export
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.c2                 (),                                               //           (terminated)
		.c3                 (),                                               //           (terminated)
		.c4                 (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	elimax_ghrd_nios_sys_clear clear (
		.clk        (clock_bridge_0_out_clk_clk),            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_clear_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_clear_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_clear_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_clear_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_clear_s1_readdata),   //                    .readdata
		.out_port   (clear_external_connection_export)       // external_connection.export
	);

	elimax_ghrd_nios_sys_jtag_uart_0 jtag_uart_0 (
		.clk            (clock_bridge_0_out_clk_clk),                                  //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	elimax_ghrd_nios_sys_led led (
		.clk        (clock_bridge_0_out_clk_clk),          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	elimax_ghrd_nios_sys_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clock_bridge_0_out_clk_clk),                                 //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	elimax_ghrd_nios_sys_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clock_bridge_0_out_clk_clk),                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	opencores_i2c opencores_i2c_0 (
		.wb_clk_i   (clock_bridge_0_out_clk_clk),                                   //            clock.clk
		.wb_rst_i   (rst_controller_001_reset_out_reset),                           //      clock_reset.reset
		.scl_pad_io (opencores_i2c_0_export_0_scl_pad_io),                          //         export_0.export
		.sda_pad_io (opencores_i2c_0_export_0_sda_pad_io),                          //                 .export
		.wb_adr_i   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver0_irq)                                      // interrupt_sender.irq
	);

	elimax_ghrd_nios_sys_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clock_bridge_0_out_clk_clk),                            //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	elimax_ghrd_nios_sys_trigger trigger (
		.clk        (clock_bridge_0_out_clk_clk),              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_trigger_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_trigger_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_trigger_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_trigger_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_trigger_s1_readdata),   //                    .readdata
		.out_port   (trigger_external_connection_export)       // external_connection.export
	);

	usb_streaming usb_streaming_0 (
		.stream_data  (usb_streaming_0_asi_in0_data),          //    asi_in0.data
		.stream_eop   (usb_streaming_0_asi_in0_endofpacket),   //           .endofpacket
		.stream_sop   (usb_streaming_0_asi_in0_startofpacket), //           .startofpacket
		.stream_valid (usb_streaming_0_asi_in0_valid),         //           .valid
		.clk          (clock_bridge_0_out_clk_clk),            //      clock.clk
		.reset_n      (~rst_controller_001_reset_out_reset),   //      reset.reset_n
		.ctl0         (usb_streaming_0_ctl0_conduit),          //       ctl0.conduit
		.clear_fifo   (usb_streaming_0_clear_fifo_conduit),    // clear_fifo.conduit
		.ctl1         (usb_streaming_0_ctl1_conduit),          //       ctl1.conduit
		.ctl2         (usb_streaming_0_ctl2_conduit),          //       ctl2.conduit
		.ctl3         (usb_streaming_0_ctl3_conduit),          //       ctl3.conduit
		.ctl5         (usb_streaming_0_ctl5_conduit),          //       ctl5.conduit
		.ctl6         (usb_streaming_0_ctl6_conduit),          //       ctl6.conduit
		.ctl7         (usb_streaming_0_ctl7_conduit),          //       ctl7.conduit
		.ctl8         (usb_streaming_0_ctl8_conduit),          //       ctl8.conduit
		.ctl11        (usb_streaming_0_ctl11_conduit),         //      ctl11.conduit
		.ctl12        (usb_streaming_0_ctl12_conduit),         //      ctl12.conduit
		.usb_data     (usb_streaming_0_usb_data_conduit),      //   usb_data.conduit
		.ctl4_sw      (usb_streaming_0_ctl4_sw_conduit)        //    ctl4_sw.conduit
	);

	elimax_ghrd_nios_sys_usbstatus usbstatus (
		.clk        (clock_bridge_0_out_clk_clk),                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_usbstatus_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_usbstatus_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_usbstatus_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_usbstatus_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_usbstatus_s1_readdata),   //                    .readdata
		.in_port    (usbstatus_external_connection_export)       // external_connection.export
	);

	videosampler #(
		.DATA_WIDTH         (32),
		.PIXEL_WIDTH        (8),
		.FIFO_DEPTH         (2048),
		.DEFAULT_SCR        (0),
		.DEFAULT_FLOWLENGTH (262144),
		.HREF_POLARITY      ("high"),
		.VSYNC_POLARITY     ("high")
	) videosampler_0 (
		.addr_rel_i (mm_interconnect_0_videosampler_0_avalon_slave_0_address),   //          avalon_slave_0.address
		.wr_i       (mm_interconnect_0_videosampler_0_avalon_slave_0_write),     //                        .write
		.datawr_i   (mm_interconnect_0_videosampler_0_avalon_slave_0_writedata), //                        .writedata
		.rd_i       (mm_interconnect_0_videosampler_0_avalon_slave_0_read),      //                        .read
		.datard_o   (mm_interconnect_0_videosampler_0_avalon_slave_0_readdata),  //                        .readdata
		.clk_i      (clock_bridge_0_out_clk_clk),                                //              clock_sink.clk
		.reset_n_i  (~rst_controller_001_reset_out_reset),                       //              reset_sink.reset_n
		.pixel_i    (videosampler_0_pixel_i_conduit),                            //                 pixel_i.conduit
		.vsync_i    (videosampler_0_vsync_i_conduit),                            //                 vsync_i.conduit
		.pclk_i     (videosampler_0_pclk_i_conduit),                             //                  pclk_i.conduit
		.href_i     (videosampler_0_href_conduit),                               //                    href.conduit
		.out_data   (videosampler_0_avalon_streaming_source_data),               // avalon_streaming_source.data
		.out_dv     (videosampler_0_avalon_streaming_source_valid),              //                        .valid
		.out_eop    (videosampler_0_avalon_streaming_source_endofpacket),        //                        .endofpacket
		.out_sop    (videosampler_0_avalon_streaming_source_startofpacket)       //                        .startofpacket
	);

	elimax_ghrd_nios_sys_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c1_clk                                            (clock_bridge_0_out_clk_clk),                                    //                                          altpll_0_c1.clk
		.clk_0_clk_clk                                              (clk_clk),                                                       //                                            clk_0_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.jtag_uart_0_reset_reset_bridge_in_reset_reset              (rst_controller_001_reset_out_reset),                            //              jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset             (rst_controller_002_reset_out_reset),                            //             nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                           (nios2_gen2_0_data_master_address),                              //                             nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                          //                                                     .waitrequest
		.nios2_gen2_0_data_master_byteenable                        (nios2_gen2_0_data_master_byteenable),                           //                                                     .byteenable
		.nios2_gen2_0_data_master_read                              (nios2_gen2_0_data_master_read),                                 //                                                     .read
		.nios2_gen2_0_data_master_readdata                          (nios2_gen2_0_data_master_readdata),                             //                                                     .readdata
		.nios2_gen2_0_data_master_write                             (nios2_gen2_0_data_master_write),                                //                                                     .write
		.nios2_gen2_0_data_master_writedata                         (nios2_gen2_0_data_master_writedata),                            //                                                     .writedata
		.nios2_gen2_0_data_master_debugaccess                       (nios2_gen2_0_data_master_debugaccess),                          //                                                     .debugaccess
		.nios2_gen2_0_instruction_master_address                    (nios2_gen2_0_instruction_master_address),                       //                      nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                (nios2_gen2_0_instruction_master_waitrequest),                   //                                                     .waitrequest
		.nios2_gen2_0_instruction_master_read                       (nios2_gen2_0_instruction_master_read),                          //                                                     .read
		.nios2_gen2_0_instruction_master_readdata                   (nios2_gen2_0_instruction_master_readdata),                      //                                                     .readdata
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),                  //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                    //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                     //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),                 //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),                //                                                     .writedata
		.clear_s1_address                                           (mm_interconnect_0_clear_s1_address),                            //                                             clear_s1.address
		.clear_s1_write                                             (mm_interconnect_0_clear_s1_write),                              //                                                     .write
		.clear_s1_readdata                                          (mm_interconnect_0_clear_s1_readdata),                           //                                                     .readdata
		.clear_s1_writedata                                         (mm_interconnect_0_clear_s1_writedata),                          //                                                     .writedata
		.clear_s1_chipselect                                        (mm_interconnect_0_clear_s1_chipselect),                         //                                                     .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),       //                        jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),         //                                                     .write
		.jtag_uart_0_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),          //                                                     .read
		.jtag_uart_0_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),      //                                                     .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),     //                                                     .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),   //                                                     .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),    //                                                     .chipselect
		.led_s1_address                                             (mm_interconnect_0_led_s1_address),                              //                                               led_s1.address
		.led_s1_write                                               (mm_interconnect_0_led_s1_write),                                //                                                     .write
		.led_s1_readdata                                            (mm_interconnect_0_led_s1_readdata),                             //                                                     .readdata
		.led_s1_writedata                                           (mm_interconnect_0_led_s1_writedata),                            //                                                     .writedata
		.led_s1_chipselect                                          (mm_interconnect_0_led_s1_chipselect),                           //                                                     .chipselect
		.nios2_gen2_0_debug_mem_slave_address                       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),        //                         nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),          //                                                     .write
		.nios2_gen2_0_debug_mem_slave_read                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),           //                                                     .read
		.nios2_gen2_0_debug_mem_slave_readdata                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),       //                                                     .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),      //                                                     .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),     //                                                     .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),    //                                                     .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),    //                                                     .debugaccess
		.onchip_memory2_0_s1_address                                (mm_interconnect_0_onchip_memory2_0_s1_address),                 //                                  onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                  (mm_interconnect_0_onchip_memory2_0_s1_write),                   //                                                     .write
		.onchip_memory2_0_s1_readdata                               (mm_interconnect_0_onchip_memory2_0_s1_readdata),                //                                                     .readdata
		.onchip_memory2_0_s1_writedata                              (mm_interconnect_0_onchip_memory2_0_s1_writedata),               //                                                     .writedata
		.onchip_memory2_0_s1_byteenable                             (mm_interconnect_0_onchip_memory2_0_s1_byteenable),              //                                                     .byteenable
		.onchip_memory2_0_s1_chipselect                             (mm_interconnect_0_onchip_memory2_0_s1_chipselect),              //                                                     .chipselect
		.onchip_memory2_0_s1_clken                                  (mm_interconnect_0_onchip_memory2_0_s1_clken),                   //                                                     .clken
		.opencores_i2c_0_avalon_slave_0_address                     (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address),      //                       opencores_i2c_0_avalon_slave_0.address
		.opencores_i2c_0_avalon_slave_0_write                       (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write),        //                                                     .write
		.opencores_i2c_0_avalon_slave_0_readdata                    (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata),     //                                                     .readdata
		.opencores_i2c_0_avalon_slave_0_writedata                   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata),    //                                                     .writedata
		.opencores_i2c_0_avalon_slave_0_waitrequest                 (~mm_interconnect_0_opencores_i2c_0_avalon_slave_0_waitrequest), //                                                     .waitrequest
		.opencores_i2c_0_avalon_slave_0_chipselect                  (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect),   //                                                     .chipselect
		.sysid_qsys_0_control_slave_address                         (mm_interconnect_0_sysid_qsys_0_control_slave_address),          //                           sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                        (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),         //                                                     .readdata
		.trigger_s1_address                                         (mm_interconnect_0_trigger_s1_address),                          //                                           trigger_s1.address
		.trigger_s1_write                                           (mm_interconnect_0_trigger_s1_write),                            //                                                     .write
		.trigger_s1_readdata                                        (mm_interconnect_0_trigger_s1_readdata),                         //                                                     .readdata
		.trigger_s1_writedata                                       (mm_interconnect_0_trigger_s1_writedata),                        //                                                     .writedata
		.trigger_s1_chipselect                                      (mm_interconnect_0_trigger_s1_chipselect),                       //                                                     .chipselect
		.usbstatus_s1_address                                       (mm_interconnect_0_usbstatus_s1_address),                        //                                         usbstatus_s1.address
		.usbstatus_s1_write                                         (mm_interconnect_0_usbstatus_s1_write),                          //                                                     .write
		.usbstatus_s1_readdata                                      (mm_interconnect_0_usbstatus_s1_readdata),                       //                                                     .readdata
		.usbstatus_s1_writedata                                     (mm_interconnect_0_usbstatus_s1_writedata),                      //                                                     .writedata
		.usbstatus_s1_chipselect                                    (mm_interconnect_0_usbstatus_s1_chipselect),                     //                                                     .chipselect
		.videosampler_0_avalon_slave_0_address                      (mm_interconnect_0_videosampler_0_avalon_slave_0_address),       //                        videosampler_0_avalon_slave_0.address
		.videosampler_0_avalon_slave_0_write                        (mm_interconnect_0_videosampler_0_avalon_slave_0_write),         //                                                     .write
		.videosampler_0_avalon_slave_0_read                         (mm_interconnect_0_videosampler_0_avalon_slave_0_read),          //                                                     .read
		.videosampler_0_avalon_slave_0_readdata                     (mm_interconnect_0_videosampler_0_avalon_slave_0_readdata),      //                                                     .readdata
		.videosampler_0_avalon_slave_0_writedata                    (mm_interconnect_0_videosampler_0_avalon_slave_0_writedata)      //                                                     .writedata
	);

	elimax_ghrd_nios_sys_irq_mapper irq_mapper (
		.clk           (clock_bridge_0_out_clk_clk),         //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clock_bridge_0_out_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clock_bridge_0_out_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
