-- elimax_ghrd_nios_sys.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity elimax_ghrd_nios_sys is
	port (
		altpll_0_areset_conduit_export       : in    std_logic                     := '0';             --       altpll_0_areset_conduit.export
		altpll_0_c0_clk                      : out   std_logic;                                        --                   altpll_0_c0.clk
		altpll_0_locked_conduit_export       : out   std_logic;                                        --       altpll_0_locked_conduit.export
		clear_external_connection_export     : out   std_logic;                                        --     clear_external_connection.export
		clk_clk                              : in    std_logic                     := '0';             --                           clk.clk
		clock_bridge_0_out_clk_clk           : out   std_logic;                                        --        clock_bridge_0_out_clk.clk
		led_external_connection_export       : out   std_logic_vector(1 downto 0);                     --       led_external_connection.export
		opencores_i2c_0_export_0_scl_pad_io  : inout std_logic                     := '0';             --      opencores_i2c_0_export_0.scl_pad_io
		opencores_i2c_0_export_0_sda_pad_io  : inout std_logic                     := '0';             --                              .sda_pad_io
		reset_reset_n                        : in    std_logic                     := '0';             --                         reset.reset_n
		trigger_external_connection_export   : out   std_logic;                                        --   trigger_external_connection.export
		usb_streaming_0_clear_fifo_conduit   : in    std_logic                     := '0';             --    usb_streaming_0_clear_fifo.conduit
		usb_streaming_0_ctl0_conduit         : out   std_logic;                                        --          usb_streaming_0_ctl0.conduit
		usb_streaming_0_ctl1_conduit         : out   std_logic;                                        --          usb_streaming_0_ctl1.conduit
		usb_streaming_0_ctl11_conduit        : out   std_logic;                                        --         usb_streaming_0_ctl11.conduit
		usb_streaming_0_ctl12_conduit        : out   std_logic;                                        --         usb_streaming_0_ctl12.conduit
		usb_streaming_0_ctl2_conduit         : out   std_logic;                                        --          usb_streaming_0_ctl2.conduit
		usb_streaming_0_ctl3_conduit         : out   std_logic;                                        --          usb_streaming_0_ctl3.conduit
		usb_streaming_0_ctl4_sw_conduit      : in    std_logic                     := '0';             --       usb_streaming_0_ctl4_sw.conduit
		usb_streaming_0_ctl5_conduit         : in    std_logic                     := '0';             --          usb_streaming_0_ctl5.conduit
		usb_streaming_0_ctl6_conduit         : in    std_logic                     := '0';             --          usb_streaming_0_ctl6.conduit
		usb_streaming_0_ctl7_conduit         : out   std_logic;                                        --          usb_streaming_0_ctl7.conduit
		usb_streaming_0_ctl8_conduit         : in    std_logic                     := '0';             --          usb_streaming_0_ctl8.conduit
		usb_streaming_0_usb_data_conduit     : inout std_logic_vector(15 downto 0) := (others => '0'); --      usb_streaming_0_usb_data.conduit
		usbstatus_external_connection_export : in    std_logic_vector(3 downto 0)  := (others => '0'); -- usbstatus_external_connection.export
		videosampler_0_href_conduit          : in    std_logic                     := '0';             --           videosampler_0_href.conduit
		videosampler_0_pclk_i_conduit        : in    std_logic                     := '0';             --         videosampler_0_pclk_i.conduit
		videosampler_0_pixel_i_conduit       : in    std_logic_vector(7 downto 0)  := (others => '0'); --        videosampler_0_pixel_i.conduit
		videosampler_0_vsync_i_conduit       : in    std_logic                     := '0'              --        videosampler_0_vsync_i.conduit
	);
end entity elimax_ghrd_nios_sys;

architecture rtl of elimax_ghrd_nios_sys is
	component IP_Filtre_Moyenneur is
		port (
			in_data    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			in_dv      : in  std_logic                     := 'X';             -- valid
			in_sop     : in  std_logic                     := 'X';             -- startofpacket
			in_eop     : in  std_logic                     := 'X';             -- endofpacket
			out_data   : out std_logic_vector(7 downto 0);                     -- data
			out_dv     : out std_logic;                                        -- valid
			out_eop    : out std_logic;                                        -- endofpacket
			out_sop    : out std_logic;                                        -- startofpacket
			CLOCK      : in  std_logic                     := 'X';             -- clk
			RESET_N    : in  std_logic                     := 'X';             -- reset_n
			addr       : in  std_logic                     := 'X';             -- address
			write_data : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read_data  : out std_logic_vector(31 downto 0);                    -- readdata
			a_read     : in  std_logic                     := 'X';             -- read
			a_write    : in  std_logic                     := 'X'              -- write
		);
	end component IP_Filtre_Moyenneur;

	component elimax_ghrd_nios_sys_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component elimax_ghrd_nios_sys_altpll_0;

	component elimax_ghrd_nios_sys_clear is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component elimax_ghrd_nios_sys_clear;

	component elimax_ghrd_nios_sys_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component elimax_ghrd_nios_sys_jtag_uart_0;

	component elimax_ghrd_nios_sys_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(1 downto 0)                      -- export
		);
	end component elimax_ghrd_nios_sys_led;

	component elimax_ghrd_nios_sys_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(18 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(18 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component elimax_ghrd_nios_sys_nios2_gen2_0;

	component elimax_ghrd_nios_sys_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component elimax_ghrd_nios_sys_onchip_memory2_0;

	component opencores_i2c is
		port (
			wb_clk_i   : in    std_logic                    := 'X';             -- clk
			wb_rst_i   : in    std_logic                    := 'X';             -- reset
			scl_pad_io : inout std_logic                    := 'X';             -- export
			sda_pad_io : inout std_logic                    := 'X';             -- export
			wb_adr_i   : in    std_logic_vector(2 downto 0) := (others => 'X'); -- address
			wb_dat_i   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			wb_dat_o   : out   std_logic_vector(7 downto 0);                    -- readdata
			wb_we_i    : in    std_logic                    := 'X';             -- write
			wb_stb_i   : in    std_logic                    := 'X';             -- chipselect
			wb_ack_o   : out   std_logic;                                       -- waitrequest_n
			wb_inta_o  : out   std_logic                                        -- irq
		);
	end component opencores_i2c;

	component elimax_ghrd_nios_sys_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component elimax_ghrd_nios_sys_sysid_qsys_0;

	component elimax_ghrd_nios_sys_trigger is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component elimax_ghrd_nios_sys_trigger;

	component usb_streaming is
		port (
			stream_data  : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			stream_eop   : in    std_logic                     := 'X';             -- endofpacket
			stream_sop   : in    std_logic                     := 'X';             -- startofpacket
			stream_valid : in    std_logic                     := 'X';             -- valid
			clk          : in    std_logic                     := 'X';             -- clk
			reset_n      : in    std_logic                     := 'X';             -- reset_n
			ctl0         : out   std_logic;                                        -- conduit
			clear_fifo   : in    std_logic                     := 'X';             -- conduit
			ctl1         : out   std_logic;                                        -- conduit
			ctl2         : out   std_logic;                                        -- conduit
			ctl3         : out   std_logic;                                        -- conduit
			ctl5         : in    std_logic                     := 'X';             -- conduit
			ctl6         : in    std_logic                     := 'X';             -- conduit
			ctl7         : out   std_logic;                                        -- conduit
			ctl8         : in    std_logic                     := 'X';             -- conduit
			ctl11        : out   std_logic;                                        -- conduit
			ctl12        : out   std_logic;                                        -- conduit
			usb_data     : inout std_logic_vector(15 downto 0) := (others => 'X'); -- conduit
			ctl4_sw      : in    std_logic                     := 'X'              -- conduit
		);
	end component usb_streaming;

	component elimax_ghrd_nios_sys_usbstatus is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component elimax_ghrd_nios_sys_usbstatus;

	component videosampler is
		generic (
			DATA_WIDTH         : integer := 32;
			PIXEL_WIDTH        : integer := 8;
			FIFO_DEPTH         : integer := 2048;
			DEFAULT_SCR        : integer := 0;
			DEFAULT_FLOWLENGTH : integer := 262144;
			HREF_POLARITY      : string  := "high";
			VSYNC_POLARITY     : string  := "high"
		);
		port (
			addr_rel_i : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wr_i       : in  std_logic                     := 'X';             -- write
			datawr_i   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			rd_i       : in  std_logic                     := 'X';             -- read
			datard_o   : out std_logic_vector(31 downto 0);                    -- readdata
			clk_i      : in  std_logic                     := 'X';             -- clk
			reset_n_i  : in  std_logic                     := 'X';             -- reset_n
			pixel_i    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- conduit
			vsync_i    : in  std_logic                     := 'X';             -- conduit
			pclk_i     : in  std_logic                     := 'X';             -- conduit
			href_i     : in  std_logic                     := 'X';             -- conduit
			out_data   : out std_logic_vector(7 downto 0);                     -- data
			out_dv     : out std_logic;                                        -- valid
			out_eop    : out std_logic;                                        -- endofpacket
			out_sop    : out std_logic                                         -- startofpacket
		);
	end component videosampler;

	component elimax_ghrd_nios_sys_mm_interconnect_0 is
		port (
			altpll_0_c1_clk                                            : in  std_logic                     := 'X';             -- clk
			clk_0_clk_clk                                              : in  std_logic                     := 'X';             -- clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset              : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                           : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                       : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                              : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                             : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                       : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                    : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest                : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                       : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			altpll_0_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			altpll_0_pll_slave_write                                   : out std_logic;                                        -- write
			altpll_0_pll_slave_read                                    : out std_logic;                                        -- read
			altpll_0_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_0_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			clear_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			clear_s1_write                                             : out std_logic;                                        -- write
			clear_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			clear_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			clear_s1_chipselect                                        : out std_logic;                                        -- chipselect
			IP_custom_0_avalon_slave_0_address                         : out std_logic_vector(0 downto 0);                     -- address
			IP_custom_0_avalon_slave_0_write                           : out std_logic;                                        -- write
			IP_custom_0_avalon_slave_0_read                            : out std_logic;                                        -- read
			IP_custom_0_avalon_slave_0_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			IP_custom_0_avalon_slave_0_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_address                      : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                        : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                         : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                   : out std_logic;                                        -- chipselect
			led_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			led_s1_write                                               : out std_logic;                                        -- write
			led_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_s1_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			led_s1_chipselect                                          : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                       : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                         : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                          : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                    : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                   : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                                : out std_logic_vector(14 downto 0);                    -- address
			onchip_memory2_0_s1_write                                  : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                             : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                                  : out std_logic;                                        -- clken
			opencores_i2c_0_avalon_slave_0_address                     : out std_logic_vector(2 downto 0);                     -- address
			opencores_i2c_0_avalon_slave_0_write                       : out std_logic;                                        -- write
			opencores_i2c_0_avalon_slave_0_readdata                    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			opencores_i2c_0_avalon_slave_0_writedata                   : out std_logic_vector(7 downto 0);                     -- writedata
			opencores_i2c_0_avalon_slave_0_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			opencores_i2c_0_avalon_slave_0_chipselect                  : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address                         : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			trigger_s1_address                                         : out std_logic_vector(2 downto 0);                     -- address
			trigger_s1_write                                           : out std_logic;                                        -- write
			trigger_s1_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			trigger_s1_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			trigger_s1_chipselect                                      : out std_logic;                                        -- chipselect
			usbstatus_s1_address                                       : out std_logic_vector(1 downto 0);                     -- address
			usbstatus_s1_write                                         : out std_logic;                                        -- write
			usbstatus_s1_readdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			usbstatus_s1_writedata                                     : out std_logic_vector(31 downto 0);                    -- writedata
			usbstatus_s1_chipselect                                    : out std_logic;                                        -- chipselect
			videosampler_0_avalon_slave_0_address                      : out std_logic_vector(2 downto 0);                     -- address
			videosampler_0_avalon_slave_0_write                        : out std_logic;                                        -- write
			videosampler_0_avalon_slave_0_read                         : out std_logic;                                        -- read
			videosampler_0_avalon_slave_0_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			videosampler_0_avalon_slave_0_writedata                    : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component elimax_ghrd_nios_sys_mm_interconnect_0;

	component elimax_ghrd_nios_sys_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component elimax_ghrd_nios_sys_irq_mapper;

	component elimax_ghrd_nios_sys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component elimax_ghrd_nios_sys_rst_controller;

	component elimax_ghrd_nios_sys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component elimax_ghrd_nios_sys_rst_controller_001;

	component elimax_ghrd_nios_sys_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component elimax_ghrd_nios_sys_rst_controller_002;

	signal ip_custom_0_avalon_streaming_source_valid                       : std_logic;                     -- IP_custom_0:out_dv -> usb_streaming_0:stream_valid
	signal ip_custom_0_avalon_streaming_source_data                        : std_logic_vector(7 downto 0);  -- IP_custom_0:out_data -> usb_streaming_0:stream_data
	signal ip_custom_0_avalon_streaming_source_startofpacket               : std_logic;                     -- IP_custom_0:out_sop -> usb_streaming_0:stream_sop
	signal ip_custom_0_avalon_streaming_source_endofpacket                 : std_logic;                     -- IP_custom_0:out_eop -> usb_streaming_0:stream_eop
	signal videosampler_0_avalon_streaming_source_valid                    : std_logic;                     -- videosampler_0:out_dv -> IP_custom_0:in_dv
	signal videosampler_0_avalon_streaming_source_data                     : std_logic_vector(7 downto 0);  -- videosampler_0:out_data -> IP_custom_0:in_data
	signal videosampler_0_avalon_streaming_source_startofpacket            : std_logic;                     -- videosampler_0:out_sop -> IP_custom_0:in_sop
	signal videosampler_0_avalon_streaming_source_endofpacket              : std_logic;                     -- videosampler_0:out_eop -> IP_custom_0:in_eop
	signal altpll_0_c1_clk                                                 : std_logic;                     -- altpll_0:c1 -> [clock_bridge_0_out_clk_clk, IP_custom_0:CLOCK, clear:clk, irq_mapper:clk, jtag_uart_0:clk, led:clk, mm_interconnect_0:altpll_0_c1_clk, nios2_gen2_0:clk, onchip_memory2_0:clk, opencores_i2c_0:wb_clk_i, rst_controller:clk, rst_controller_002:clk, sysid_qsys_0:clock, trigger:clk, usb_streaming_0:clk, usbstatus:clk, videosampler_0:clk_i]
	signal nios2_gen2_0_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                            : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                : std_logic_vector(18 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                   : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                  : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                              : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                         : std_logic_vector(18 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                            : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect     : std_logic;                     -- mm_interconnect_0:opencores_i2c_0_avalon_slave_0_chipselect -> opencores_i2c_0:wb_stb_i
	signal mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata       : std_logic_vector(7 downto 0);  -- opencores_i2c_0:wb_dat_o -> mm_interconnect_0:opencores_i2c_0_avalon_slave_0_readdata
	signal opencores_i2c_0_avalon_slave_0_waitrequest                      : std_logic;                     -- opencores_i2c_0:wb_ack_o -> opencores_i2c_0_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:opencores_i2c_0_avalon_slave_0_address -> opencores_i2c_0:wb_adr_i
	signal mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write          : std_logic;                     -- mm_interconnect_0:opencores_i2c_0_avalon_slave_0_write -> opencores_i2c_0:wb_we_i
	signal mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata      : std_logic_vector(7 downto 0);  -- mm_interconnect_0:opencores_i2c_0_avalon_slave_0_writedata -> opencores_i2c_0:wb_dat_i
	signal mm_interconnect_0_videosampler_0_avalon_slave_0_readdata        : std_logic_vector(31 downto 0); -- videosampler_0:datard_o -> mm_interconnect_0:videosampler_0_avalon_slave_0_readdata
	signal mm_interconnect_0_videosampler_0_avalon_slave_0_address         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:videosampler_0_avalon_slave_0_address -> videosampler_0:addr_rel_i
	signal mm_interconnect_0_videosampler_0_avalon_slave_0_read            : std_logic;                     -- mm_interconnect_0:videosampler_0_avalon_slave_0_read -> videosampler_0:rd_i
	signal mm_interconnect_0_videosampler_0_avalon_slave_0_write           : std_logic;                     -- mm_interconnect_0:videosampler_0_avalon_slave_0_write -> videosampler_0:wr_i
	signal mm_interconnect_0_videosampler_0_avalon_slave_0_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:videosampler_0_avalon_slave_0_writedata -> videosampler_0:datawr_i
	signal mm_interconnect_0_ip_custom_0_avalon_slave_0_readdata           : std_logic_vector(31 downto 0); -- IP_custom_0:read_data -> mm_interconnect_0:IP_custom_0_avalon_slave_0_readdata
	signal mm_interconnect_0_ip_custom_0_avalon_slave_0_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:IP_custom_0_avalon_slave_0_address -> IP_custom_0:addr
	signal mm_interconnect_0_ip_custom_0_avalon_slave_0_read               : std_logic;                     -- mm_interconnect_0:IP_custom_0_avalon_slave_0_read -> IP_custom_0:a_read
	signal mm_interconnect_0_ip_custom_0_avalon_slave_0_write              : std_logic;                     -- mm_interconnect_0:IP_custom_0_avalon_slave_0_write -> IP_custom_0:a_write
	signal mm_interconnect_0_ip_custom_0_avalon_slave_0_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:IP_custom_0_avalon_slave_0_writedata -> IP_custom_0:write_data
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata           : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest      : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_altpll_0_pll_slave_readdata                   : std_logic_vector(31 downto 0); -- altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	signal mm_interconnect_0_altpll_0_pll_slave_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	signal mm_interconnect_0_altpll_0_pll_slave_read                       : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	signal mm_interconnect_0_altpll_0_pll_slave_write                      : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	signal mm_interconnect_0_altpll_0_pll_slave_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                  : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                   : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_trigger_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:trigger_s1_chipselect -> trigger:chipselect
	signal mm_interconnect_0_trigger_s1_readdata                           : std_logic_vector(31 downto 0); -- trigger:readdata -> mm_interconnect_0:trigger_s1_readdata
	signal mm_interconnect_0_trigger_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:trigger_s1_address -> trigger:address
	signal mm_interconnect_0_trigger_s1_write                              : std_logic;                     -- mm_interconnect_0:trigger_s1_write -> mm_interconnect_0_trigger_s1_write:in
	signal mm_interconnect_0_trigger_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:trigger_s1_writedata -> trigger:writedata
	signal mm_interconnect_0_clear_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:clear_s1_chipselect -> clear:chipselect
	signal mm_interconnect_0_clear_s1_readdata                             : std_logic_vector(31 downto 0); -- clear:readdata -> mm_interconnect_0:clear_s1_readdata
	signal mm_interconnect_0_clear_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:clear_s1_address -> clear:address
	signal mm_interconnect_0_clear_s1_write                                : std_logic;                     -- mm_interconnect_0:clear_s1_write -> mm_interconnect_0_clear_s1_write:in
	signal mm_interconnect_0_clear_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:clear_s1_writedata -> clear:writedata
	signal mm_interconnect_0_led_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:led_s1_chipselect -> led:chipselect
	signal mm_interconnect_0_led_s1_readdata                               : std_logic_vector(31 downto 0); -- led:readdata -> mm_interconnect_0:led_s1_readdata
	signal mm_interconnect_0_led_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_s1_address -> led:address
	signal mm_interconnect_0_led_s1_write                                  : std_logic;                     -- mm_interconnect_0:led_s1_write -> mm_interconnect_0_led_s1_write:in
	signal mm_interconnect_0_led_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_s1_writedata -> led:writedata
	signal mm_interconnect_0_usbstatus_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:usbstatus_s1_chipselect -> usbstatus:chipselect
	signal mm_interconnect_0_usbstatus_s1_readdata                         : std_logic_vector(31 downto 0); -- usbstatus:readdata -> mm_interconnect_0:usbstatus_s1_readdata
	signal mm_interconnect_0_usbstatus_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:usbstatus_s1_address -> usbstatus:address
	signal mm_interconnect_0_usbstatus_s1_write                            : std_logic;                     -- mm_interconnect_0:usbstatus_s1_write -> mm_interconnect_0_usbstatus_s1_write:in
	signal mm_interconnect_0_usbstatus_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:usbstatus_s1_writedata -> usbstatus:writedata
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- opencores_i2c_0:wb_inta_o -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	signal nios2_gen2_0_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, opencores_i2c_0:wb_rst_i, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal rst_controller_002_reset_out_reset                              : std_logic;                     -- rst_controller_002:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset_req                          : std_logic;                     -- rst_controller_002:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]
	signal nios2_gen2_0_debug_reset_request_reset                          : std_logic;                     -- nios2_gen2_0:debug_reset_request -> rst_controller_002:reset_in1
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_opencores_i2c_0_avalon_slave_0_inv            : std_logic;                     -- opencores_i2c_0_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:opencores_i2c_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_trigger_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_trigger_s1_write:inv -> trigger:write_n
	signal mm_interconnect_0_clear_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_clear_s1_write:inv -> clear:write_n
	signal mm_interconnect_0_led_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_led_s1_write:inv -> led:write_n
	signal mm_interconnect_0_usbstatus_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_usbstatus_s1_write:inv -> usbstatus:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [IP_custom_0:RESET_N, clear:reset_n, jtag_uart_0:rst_n, led:reset_n, sysid_qsys_0:reset_n, trigger:reset_n, usb_streaming_0:reset_n, usbstatus:reset_n, videosampler_0:reset_n_i]
	signal rst_controller_002_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> nios2_gen2_0:reset_n

begin

	ip_custom_0 : component IP_Filtre_Moyenneur
		port map (
			in_data    => videosampler_0_avalon_streaming_source_data,             --   avalon_streaming_sink.data
			in_dv      => videosampler_0_avalon_streaming_source_valid,            --                        .valid
			in_sop     => videosampler_0_avalon_streaming_source_startofpacket,    --                        .startofpacket
			in_eop     => videosampler_0_avalon_streaming_source_endofpacket,      --                        .endofpacket
			out_data   => ip_custom_0_avalon_streaming_source_data,                -- avalon_streaming_source.data
			out_dv     => ip_custom_0_avalon_streaming_source_valid,               --                        .valid
			out_eop    => ip_custom_0_avalon_streaming_source_endofpacket,         --                        .endofpacket
			out_sop    => ip_custom_0_avalon_streaming_source_startofpacket,       --                        .startofpacket
			CLOCK      => altpll_0_c1_clk,                                         --              clock_sink.clk
			RESET_N    => rst_controller_reset_out_reset_ports_inv,                --              reset_sink.reset_n
			addr       => mm_interconnect_0_ip_custom_0_avalon_slave_0_address(0), --          avalon_slave_0.address
			write_data => mm_interconnect_0_ip_custom_0_avalon_slave_0_writedata,  --                        .writedata
			read_data  => mm_interconnect_0_ip_custom_0_avalon_slave_0_readdata,   --                        .readdata
			a_read     => mm_interconnect_0_ip_custom_0_avalon_slave_0_read,       --                        .read
			a_write    => mm_interconnect_0_ip_custom_0_avalon_slave_0_write       --                        .write
		);

	altpll_0 : component elimax_ghrd_nios_sys_altpll_0
		port map (
			clk                => clk_clk,                                        --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset,             -- inclk_interface_reset.reset
			read               => mm_interconnect_0_altpll_0_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_altpll_0_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_altpll_0_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_altpll_0_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_altpll_0_pll_slave_writedata, --                      .writedata
			c0                 => altpll_0_c0_clk,                                --                    c0.clk
			c1                 => altpll_0_c1_clk,                                --                    c1.clk
			areset             => altpll_0_areset_conduit_export,                 --        areset_conduit.export
			locked             => altpll_0_locked_conduit_export,                 --        locked_conduit.export
			scandone           => open,                                           --           (terminated)
			scandataout        => open,                                           --           (terminated)
			c2                 => open,                                           --           (terminated)
			c3                 => open,                                           --           (terminated)
			c4                 => open,                                           --           (terminated)
			phasedone          => open,                                           --           (terminated)
			phasecounterselect => "000",                                          --           (terminated)
			phaseupdown        => '0',                                            --           (terminated)
			phasestep          => '0',                                            --           (terminated)
			scanclk            => '0',                                            --           (terminated)
			scanclkena         => '0',                                            --           (terminated)
			scandata           => '0',                                            --           (terminated)
			configupdate       => '0'                                             --           (terminated)
		);

	clear : component elimax_ghrd_nios_sys_clear
		port map (
			clk        => altpll_0_c1_clk,                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_clear_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_clear_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_clear_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_clear_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_clear_s1_readdata,        --                    .readdata
			out_port   => clear_external_connection_export            -- external_connection.export
		);

	jtag_uart_0 : component elimax_ghrd_nios_sys_jtag_uart_0
		port map (
			clk            => altpll_0_c1_clk,                                                 --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                         --               irq.irq
		);

	led : component elimax_ghrd_nios_sys_led
		port map (
			clk        => altpll_0_c1_clk,                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_s1_readdata,        --                    .readdata
			out_port   => led_external_connection_export            -- external_connection.export
		);

	nios2_gen2_0 : component elimax_ghrd_nios_sys_nios2_gen2_0
		port map (
			clk                                 => altpll_0_c1_clk,                                            --                       clk.clk
			reset_n                             => rst_controller_002_reset_out_reset_ports_inv,               --                     reset.reset_n
			reset_req                           => rst_controller_002_reset_out_reset_req,                     --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component elimax_ghrd_nios_sys_onchip_memory2_0
		port map (
			clk        => altpll_0_c1_clk,                                  --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	opencores_i2c_0 : component opencores_i2c
		port map (
			wb_clk_i   => altpll_0_c1_clk,                                             --            clock.clk
			wb_rst_i   => rst_controller_reset_out_reset,                              --      clock_reset.reset
			scl_pad_io => opencores_i2c_0_export_0_scl_pad_io,                         --         export_0.export
			sda_pad_io => opencores_i2c_0_export_0_sda_pad_io,                         --                 .export
			wb_adr_i   => mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => opencores_i2c_0_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			wb_inta_o  => irq_mapper_receiver0_irq                                     -- interrupt_sender.irq
		);

	sysid_qsys_0 : component elimax_ghrd_nios_sys_sysid_qsys_0
		port map (
			clock    => altpll_0_c1_clk,                                         --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	trigger : component elimax_ghrd_nios_sys_trigger
		port map (
			clk        => altpll_0_c1_clk,                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_trigger_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_trigger_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_trigger_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_trigger_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_trigger_s1_readdata,        --                    .readdata
			out_port   => trigger_external_connection_export            -- external_connection.export
		);

	usb_streaming_0 : component usb_streaming
		port map (
			stream_data  => ip_custom_0_avalon_streaming_source_data,          --    asi_in0.data
			stream_eop   => ip_custom_0_avalon_streaming_source_endofpacket,   --           .endofpacket
			stream_sop   => ip_custom_0_avalon_streaming_source_startofpacket, --           .startofpacket
			stream_valid => ip_custom_0_avalon_streaming_source_valid,         --           .valid
			clk          => altpll_0_c1_clk,                                   --      clock.clk
			reset_n      => rst_controller_reset_out_reset_ports_inv,          --      reset.reset_n
			ctl0         => usb_streaming_0_ctl0_conduit,                      --       ctl0.conduit
			clear_fifo   => usb_streaming_0_clear_fifo_conduit,                -- clear_fifo.conduit
			ctl1         => usb_streaming_0_ctl1_conduit,                      --       ctl1.conduit
			ctl2         => usb_streaming_0_ctl2_conduit,                      --       ctl2.conduit
			ctl3         => usb_streaming_0_ctl3_conduit,                      --       ctl3.conduit
			ctl5         => usb_streaming_0_ctl5_conduit,                      --       ctl5.conduit
			ctl6         => usb_streaming_0_ctl6_conduit,                      --       ctl6.conduit
			ctl7         => usb_streaming_0_ctl7_conduit,                      --       ctl7.conduit
			ctl8         => usb_streaming_0_ctl8_conduit,                      --       ctl8.conduit
			ctl11        => usb_streaming_0_ctl11_conduit,                     --      ctl11.conduit
			ctl12        => usb_streaming_0_ctl12_conduit,                     --      ctl12.conduit
			usb_data     => usb_streaming_0_usb_data_conduit,                  --   usb_data.conduit
			ctl4_sw      => usb_streaming_0_ctl4_sw_conduit                    --    ctl4_sw.conduit
		);

	usbstatus : component elimax_ghrd_nios_sys_usbstatus
		port map (
			clk        => altpll_0_c1_clk,                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_usbstatus_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_usbstatus_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_usbstatus_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_usbstatus_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_usbstatus_s1_readdata,        --                    .readdata
			in_port    => usbstatus_external_connection_export            -- external_connection.export
		);

	videosampler_0 : component videosampler
		generic map (
			DATA_WIDTH         => 32,
			PIXEL_WIDTH        => 8,
			FIFO_DEPTH         => 2048,
			DEFAULT_SCR        => 0,
			DEFAULT_FLOWLENGTH => 262144,
			HREF_POLARITY      => "high",
			VSYNC_POLARITY     => "high"
		)
		port map (
			addr_rel_i => mm_interconnect_0_videosampler_0_avalon_slave_0_address,   --          avalon_slave_0.address
			wr_i       => mm_interconnect_0_videosampler_0_avalon_slave_0_write,     --                        .write
			datawr_i   => mm_interconnect_0_videosampler_0_avalon_slave_0_writedata, --                        .writedata
			rd_i       => mm_interconnect_0_videosampler_0_avalon_slave_0_read,      --                        .read
			datard_o   => mm_interconnect_0_videosampler_0_avalon_slave_0_readdata,  --                        .readdata
			clk_i      => altpll_0_c1_clk,                                           --              clock_sink.clk
			reset_n_i  => rst_controller_reset_out_reset_ports_inv,                  --              reset_sink.reset_n
			pixel_i    => videosampler_0_pixel_i_conduit,                            --                 pixel_i.conduit
			vsync_i    => videosampler_0_vsync_i_conduit,                            --                 vsync_i.conduit
			pclk_i     => videosampler_0_pclk_i_conduit,                             --                  pclk_i.conduit
			href_i     => videosampler_0_href_conduit,                               --                    href.conduit
			out_data   => videosampler_0_avalon_streaming_source_data,               -- avalon_streaming_source.data
			out_dv     => videosampler_0_avalon_streaming_source_valid,              --                        .valid
			out_eop    => videosampler_0_avalon_streaming_source_endofpacket,        --                        .endofpacket
			out_sop    => videosampler_0_avalon_streaming_source_startofpacket       --                        .startofpacket
		);

	mm_interconnect_0 : component elimax_ghrd_nios_sys_mm_interconnect_0
		port map (
			altpll_0_c1_clk                                            => altpll_0_c1_clk,                                             --                                          altpll_0_c1.clk
			clk_0_clk_clk                                              => clk_clk,                                                     --                                            clk_0_clk.clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                          -- altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset              => rst_controller_reset_out_reset,                              --              jtag_uart_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset             => rst_controller_002_reset_out_reset,                          --             nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                           => nios2_gen2_0_data_master_address,                            --                             nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                        --                                                     .waitrequest
			nios2_gen2_0_data_master_byteenable                        => nios2_gen2_0_data_master_byteenable,                         --                                                     .byteenable
			nios2_gen2_0_data_master_read                              => nios2_gen2_0_data_master_read,                               --                                                     .read
			nios2_gen2_0_data_master_readdata                          => nios2_gen2_0_data_master_readdata,                           --                                                     .readdata
			nios2_gen2_0_data_master_write                             => nios2_gen2_0_data_master_write,                              --                                                     .write
			nios2_gen2_0_data_master_writedata                         => nios2_gen2_0_data_master_writedata,                          --                                                     .writedata
			nios2_gen2_0_data_master_debugaccess                       => nios2_gen2_0_data_master_debugaccess,                        --                                                     .debugaccess
			nios2_gen2_0_instruction_master_address                    => nios2_gen2_0_instruction_master_address,                     --                      nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest                => nios2_gen2_0_instruction_master_waitrequest,                 --                                                     .waitrequest
			nios2_gen2_0_instruction_master_read                       => nios2_gen2_0_instruction_master_read,                        --                                                     .read
			nios2_gen2_0_instruction_master_readdata                   => nios2_gen2_0_instruction_master_readdata,                    --                                                     .readdata
			altpll_0_pll_slave_address                                 => mm_interconnect_0_altpll_0_pll_slave_address,                --                                   altpll_0_pll_slave.address
			altpll_0_pll_slave_write                                   => mm_interconnect_0_altpll_0_pll_slave_write,                  --                                                     .write
			altpll_0_pll_slave_read                                    => mm_interconnect_0_altpll_0_pll_slave_read,                   --                                                     .read
			altpll_0_pll_slave_readdata                                => mm_interconnect_0_altpll_0_pll_slave_readdata,               --                                                     .readdata
			altpll_0_pll_slave_writedata                               => mm_interconnect_0_altpll_0_pll_slave_writedata,              --                                                     .writedata
			clear_s1_address                                           => mm_interconnect_0_clear_s1_address,                          --                                             clear_s1.address
			clear_s1_write                                             => mm_interconnect_0_clear_s1_write,                            --                                                     .write
			clear_s1_readdata                                          => mm_interconnect_0_clear_s1_readdata,                         --                                                     .readdata
			clear_s1_writedata                                         => mm_interconnect_0_clear_s1_writedata,                        --                                                     .writedata
			clear_s1_chipselect                                        => mm_interconnect_0_clear_s1_chipselect,                       --                                                     .chipselect
			IP_custom_0_avalon_slave_0_address                         => mm_interconnect_0_ip_custom_0_avalon_slave_0_address,        --                           IP_custom_0_avalon_slave_0.address
			IP_custom_0_avalon_slave_0_write                           => mm_interconnect_0_ip_custom_0_avalon_slave_0_write,          --                                                     .write
			IP_custom_0_avalon_slave_0_read                            => mm_interconnect_0_ip_custom_0_avalon_slave_0_read,           --                                                     .read
			IP_custom_0_avalon_slave_0_readdata                        => mm_interconnect_0_ip_custom_0_avalon_slave_0_readdata,       --                                                     .readdata
			IP_custom_0_avalon_slave_0_writedata                       => mm_interconnect_0_ip_custom_0_avalon_slave_0_writedata,      --                                                     .writedata
			jtag_uart_0_avalon_jtag_slave_address                      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --                        jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                                     .write
			jtag_uart_0_avalon_jtag_slave_read                         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                                     .read
			jtag_uart_0_avalon_jtag_slave_readdata                     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                                     .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                                     .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                                     .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                                     .chipselect
			led_s1_address                                             => mm_interconnect_0_led_s1_address,                            --                                               led_s1.address
			led_s1_write                                               => mm_interconnect_0_led_s1_write,                              --                                                     .write
			led_s1_readdata                                            => mm_interconnect_0_led_s1_readdata,                           --                                                     .readdata
			led_s1_writedata                                           => mm_interconnect_0_led_s1_writedata,                          --                                                     .writedata
			led_s1_chipselect                                          => mm_interconnect_0_led_s1_chipselect,                         --                                                     .chipselect
			nios2_gen2_0_debug_mem_slave_address                       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,      --                         nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,        --                                                     .write
			nios2_gen2_0_debug_mem_slave_read                          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,         --                                                     .read
			nios2_gen2_0_debug_mem_slave_readdata                      => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,     --                                                     .readdata
			nios2_gen2_0_debug_mem_slave_writedata                     => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,    --                                                     .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,   --                                                     .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                   => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,  --                                                     .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                   => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,  --                                                     .debugaccess
			onchip_memory2_0_s1_address                                => mm_interconnect_0_onchip_memory2_0_s1_address,               --                                  onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                                  => mm_interconnect_0_onchip_memory2_0_s1_write,                 --                                                     .write
			onchip_memory2_0_s1_readdata                               => mm_interconnect_0_onchip_memory2_0_s1_readdata,              --                                                     .readdata
			onchip_memory2_0_s1_writedata                              => mm_interconnect_0_onchip_memory2_0_s1_writedata,             --                                                     .writedata
			onchip_memory2_0_s1_byteenable                             => mm_interconnect_0_onchip_memory2_0_s1_byteenable,            --                                                     .byteenable
			onchip_memory2_0_s1_chipselect                             => mm_interconnect_0_onchip_memory2_0_s1_chipselect,            --                                                     .chipselect
			onchip_memory2_0_s1_clken                                  => mm_interconnect_0_onchip_memory2_0_s1_clken,                 --                                                     .clken
			opencores_i2c_0_avalon_slave_0_address                     => mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address,    --                       opencores_i2c_0_avalon_slave_0.address
			opencores_i2c_0_avalon_slave_0_write                       => mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write,      --                                                     .write
			opencores_i2c_0_avalon_slave_0_readdata                    => mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata,   --                                                     .readdata
			opencores_i2c_0_avalon_slave_0_writedata                   => mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata,  --                                                     .writedata
			opencores_i2c_0_avalon_slave_0_waitrequest                 => mm_interconnect_0_opencores_i2c_0_avalon_slave_0_inv,        --                                                     .waitrequest
			opencores_i2c_0_avalon_slave_0_chipselect                  => mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect, --                                                     .chipselect
			sysid_qsys_0_control_slave_address                         => mm_interconnect_0_sysid_qsys_0_control_slave_address,        --                           sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                        => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,       --                                                     .readdata
			trigger_s1_address                                         => mm_interconnect_0_trigger_s1_address,                        --                                           trigger_s1.address
			trigger_s1_write                                           => mm_interconnect_0_trigger_s1_write,                          --                                                     .write
			trigger_s1_readdata                                        => mm_interconnect_0_trigger_s1_readdata,                       --                                                     .readdata
			trigger_s1_writedata                                       => mm_interconnect_0_trigger_s1_writedata,                      --                                                     .writedata
			trigger_s1_chipselect                                      => mm_interconnect_0_trigger_s1_chipselect,                     --                                                     .chipselect
			usbstatus_s1_address                                       => mm_interconnect_0_usbstatus_s1_address,                      --                                         usbstatus_s1.address
			usbstatus_s1_write                                         => mm_interconnect_0_usbstatus_s1_write,                        --                                                     .write
			usbstatus_s1_readdata                                      => mm_interconnect_0_usbstatus_s1_readdata,                     --                                                     .readdata
			usbstatus_s1_writedata                                     => mm_interconnect_0_usbstatus_s1_writedata,                    --                                                     .writedata
			usbstatus_s1_chipselect                                    => mm_interconnect_0_usbstatus_s1_chipselect,                   --                                                     .chipselect
			videosampler_0_avalon_slave_0_address                      => mm_interconnect_0_videosampler_0_avalon_slave_0_address,     --                        videosampler_0_avalon_slave_0.address
			videosampler_0_avalon_slave_0_write                        => mm_interconnect_0_videosampler_0_avalon_slave_0_write,       --                                                     .write
			videosampler_0_avalon_slave_0_read                         => mm_interconnect_0_videosampler_0_avalon_slave_0_read,        --                                                     .read
			videosampler_0_avalon_slave_0_readdata                     => mm_interconnect_0_videosampler_0_avalon_slave_0_readdata,    --                                                     .readdata
			videosampler_0_avalon_slave_0_writedata                    => mm_interconnect_0_videosampler_0_avalon_slave_0_writedata    --                                                     .writedata
		);

	irq_mapper : component elimax_ghrd_nios_sys_irq_mapper
		port map (
			clk           => altpll_0_c1_clk,                    --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			sender_irq    => nios2_gen2_0_irq_irq                --    sender.irq
		);

	rst_controller : component elimax_ghrd_nios_sys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => altpll_0_c1_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component elimax_ghrd_nios_sys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component elimax_ghrd_nios_sys_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => altpll_0_c1_clk,                        --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_opencores_i2c_0_avalon_slave_0_inv <= not opencores_i2c_0_avalon_slave_0_waitrequest;

	mm_interconnect_0_trigger_s1_write_ports_inv <= not mm_interconnect_0_trigger_s1_write;

	mm_interconnect_0_clear_s1_write_ports_inv <= not mm_interconnect_0_clear_s1_write;

	mm_interconnect_0_led_s1_write_ports_inv <= not mm_interconnect_0_led_s1_write;

	mm_interconnect_0_usbstatus_s1_write_ports_inv <= not mm_interconnect_0_usbstatus_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	clock_bridge_0_out_clk_clk <= altpll_0_c1_clk;

end architecture rtl; -- of elimax_ghrd_nios_sys
